`default_nettype none

module cache (
    // Global clock.
    input  wire        i_clk,
    // Synchronous active-high reset.
    input  wire        i_rst,
    // External memory interface. See hart interface for details. This
    // interface is nearly identical to the phase 5 memory interface, with the
    // exception that the byte mask (`o_mem_mask`) has been removed. This is
    // no longer needed as the cache will only access the memory at word
    // granularity, and implement masking internally.
    input  wire        i_mem_ready,
    output wire [31:0] o_mem_addr,
    output wire        o_mem_ren,
    output wire        o_mem_wen,
    output wire [31:0] o_mem_wdata,
    input  wire [31:0] i_mem_rdata,
    input  wire        i_mem_valid,

    // Interface to CPU hart. This is nearly identical to the phase 5 hart memory
    // interface, but includes a stall signal (`o_busy`), and the input/output
    // polarities are swapped for obvious reasons.
    //
    // The CPU should use this as a stall signal for both instruction fetch
    // (IF) and memory (MEM) stages, from the instruction or data cache
    // respectively. If a memory request is made (`i_req_ren` for instruction
    // cache, or either `i_req_ren` or `i_req_wen` for data cache), this
    // should be asserted *combinationally* if the request results in a cache
    // miss.
    //
    // In case of a cache miss, the CPU must stall the respective pipeline
    // stage and deassert ren/wen on subsequent cycles, until the cache
    // deasserts `o_busy` to indicate it has serviced the cache miss. However,
    // the CPU must keep the other request lines constant. For example, the
    // CPU should not change the request address while stalling.
    output wire        o_busy,
    // 32-bit read/write address to access from the cache. This should be
    // 32-bit aligned (i.e. the two LSBs should be zero). See `i_req_mask` for
    // how to perform half-word and byte accesses to unaligned addresses.
    input  wire [31:0] i_req_addr,
    // When asserted, the cache should perform a read at the aligned address
    // specified by `i_req_addr` and return the 32-bit word at that address,
    // either immediately (i.e. combinationally) on a cache hit, or
    // synchronously on a cache miss. It is illegal to assert this and
    // `i_dmem_wen` on the same cycle.
    input  wire        i_req_ren,
    // When asserted, the cache should perform a write at the aligned address
    // specified by `i_req_addr` with the 32-bit word provided in
    // `o_req_wdata` (specified by the mask). This is necessarily synchronous,
    // but may either happen on the next clock edge (on a cache hit) or after
    // multiple cycles of latency (cache miss). As the cache is write-through
    // and write-allocate, writes must be applied to both the cache and
    // underlying memory.
    // It is illegal to assert this and `i_dmem_ren` on the same cycle.
    input  wire        i_req_wen,
    // The memory interface expects word (32 bit) aligned addresses. However,
    // WISC-25 supports byte and half-word loads and stores at unaligned and
    // 16-bit aligned addresses, respectively. To support this, the access
    // mask specifies which bytes within the 32-bit word are actually read
    // from or written to memory.
    input  wire [ 3:0] i_req_mask,
    // The 32-bit word to write to memory, if the request is a write
    // (i_req_wen is asserted). Only the bytes corresponding to set bits in
    // the mask should be written into the cache (and to backing memory).
    input  wire [31:0] i_req_wdata,
    // THe 32-bit data word read from memory on a read request.
    output wire [31:0] o_res_rdata
);
  // These parameters are equivalent to those provided in the project
  // 6 specification. Feel free to use them, but hardcoding these numbers
  // rather than using the localparams is also permitted, as long as the
  // same values are used (and consistent with the project specification).
  //
  // 32 sets * 2 ways per set * 16 bytes per way = 1K cache
  localparam O = 4;  // 4 bit offset => 16 byte cache line
  localparam S = 5;  // 5 bit set index => 32 sets
  localparam DEPTH = 2 ** S;  // 32 sets
  localparam W = 2;  // 2 way set associative, NMRU
  localparam T = 32 - O - S;  // 23 bit tag
  localparam D = 2 ** O / 4;  // 16 bytes per line / 4 bytes per word = 4 words per line

  //reg versions of the outputs of the module 
  reg [31:0] o_mem_addr_reg;
  assign o_mem_addr = o_mem_addr_reg;
  reg o_mem_ren_reg;
  assign o_mem_ren = o_mem_ren_reg;
  reg o_mem_wen_reg;
  assign o_mem_wen_reg = o_mem_wen_reg;
  reg [31:0] o_mem_wdata_reg;
  assign o_mem_wdata = o_mem_wdata_reg;
  reg busy1;
  assign o_busy = busy1;

  // The following memory arrays model the cache structure. As this is
  // an internal implementation detail, you are *free* to modify these
  // arrays as you please.

  // Backing memory, modeled as two separate ways.
  reg [   31:0] datas0[DEPTH - 1:0][D - 1:0];   //stores first line in set   (32 lines x 4 words per line)
  reg [   31:0] datas1[DEPTH - 1:0][D - 1:0];  //stores second line in set 
  reg [T - 1:0] tags0[DEPTH - 1:0];  //stores tag from first line in set
  reg [T - 1:0] tags1[DEPTH - 1:0];  //stores tag from second line in set
  reg [1:0] valid [DEPTH - 1:0];  //2-bit valid (one for each line in set)
  reg       lru   [DEPTH - 1:0];  //bit to track lru

  // Fill in your implementation here.

  /*
 i_req_addr is word aligned so 2 LSBs are 0 
 */
  wire [22:0] req_tag = i_req_addr[31:9];  //top 23 bits are tag 
  wire [4:0] req_index = i_req_addr[8:4];  //5 set bits in address
  wire [1:0] req_wrdOffset = i_req_addr[3:2];  //2 bits for word offset for 16-byte blocks 
  wire hit;

  //check if valid bit is set & if tag matches request 
  wire Line0_hit = valid[req_index][0] && (tags0[req_index] == req_tag);
  wire Line1_hit = valid[req_index][1] && (tags1[req_index] == req_tag);
  assign hit = Line0_hit || Line1_hit;

  
  //FSM STATES
  localparam IDLE    = 2'b00;
  localparam MEMREAD = 2'b01;
  localparam MEMWRITE= 2'b10;
  reg [1:0] state;
  reg [1:0] next_state;

  //fsm state transition
  always @(posedge i_clk) begin
    if (i_rst) begin
      state <= IDLE;
      busy1 <= 0;
    end else begin
      state <= next_state;
    end
  end

  //Basic recap of cache organization
  //32 sets, 2 way associative with each block having 4 words
  //2 bits of the address are required to access each word, word aligned hence
  //add[3:2]
  //2 way associative implies that each set can hold 2 blocks of data
  //32 sets, hence 5 bits required to index this, or add[8:4]
  //rest of the bits are used for tag-inspection, given by [31:9]
  //
  //When a request is sent by the CPI via i_req_wen or i_req_ren, check if its
  //a hit: if hit, combinational read from the cache. 


  ///////////RESET LOGIC
  integer i, x;
  always @(posedge i_clk) begin
    if (i_rst) begin
      for (i = 0; i < 32; i = i + 1) begin
        valid[i] <= 2'd0;
        tags0[i] <= 23'd0;
        tags1[i] <= 23'd0;
        lru[i]   <= 1'd0;
        for (x = 0; x < 4; x = x + 1) begin
          datas0[i][x] <= 32'b0;
          datas1[i][x] <= 32'b0;
        end
      end
    end
  end

  reg [1:0] mem_add_read;



  //2 registers to keep track of what the request-signal type was
  reg i_req_wen_ff;
  reg i_req_ren_ff;

  //set which kind of request
  always @(posedge i_clk) begin
    if (i_rst) begin
      i_req_wen_ff <= 1'b0;
      i_req_ren_ff <= 1'b0;
    end else begin
      if (state == IDLE) begin
        i_req_wen_ff <= i_req_wen;
        i_req_ren_ff <= i_req_ren;
      end
    end
  end

  //LOGIC FOR FETCHING LINES FROM MEMORY IN MEMREAD STATE
  //if currently in the MEMREAD state, attempt to sequentially read addresses
  //for the block 
  //the data to load from memory via offset should be given by this
  wire [31:0] o_req_addr_offset;

  //cycle to include word wanted and the following three words
  assign o_req_addr_offset = i_req_addr +{28'b0, mem_add_read, 2'b0};
  

  //logic for loading 4 words of data on any read from memory
  always @(posedge i_clk) begin
    if (i_rst) begin
      mem_add_read <= 2'b0;
    end
    //if in any state other than MEMREAD, set mem_add_read to 0
    if (state != MEMREAD) begin
      mem_add_read <= 2'b0;
    end
    if (state == MEMREAD) begin
      //might need seperate state machine that goes 
      // i_mem_ready (can accept a value) -> i_mem_valid (finally fetched
      // value)-> i_mem_ready (can accept a value) etc 
      //if the current state is MEMREAD AND the value being shown by memory
      //is valid, then load it into the cache
      //increment the mem_add_read
      //
      //NOTE: is this i_mem_valid? only read the value being shown by memory
      //if its valid?
      //would i_mem_ready be false while memory is waiting/fetching?
      //if the memory is not ready maintain the current address being
      //presented to memory
      //if the memory is NOT ready for a request, maintain the current address
      //being presented to it
      if (~i_mem_ready) begin
        mem_add_read <= mem_add_read;
        o_mem_ren_reg <= 1'b0;
      end else begin 
        o_mem_addr_reg <= o_req_addr_offset;
        o_mem_ren_reg <= 1'b1;
      end
      //once memory IS ready, then present it the address. 
      //NOTE, assumes that once it reads the address, i_mem_ready goes **LOW**
      //and i_mem_valid goes **LOW**. 
      if (i_mem_valid) begin
        //TODO: logic for loading the specific word into the specific block 
        //in the cache?
        //recall that writing to a cache is sequential, hence should be in
        //a sequential block
        //uses LRU policy, so...
        //1) check if either way is empty, then allocate there
        //2) if **both** ways are not-empty, evict the LRU

        //if first line is empty
        if (~valid[req_index][0]) begin
          datas0[req_index][mem_add_read] <= i_mem_rdata;
          tags0[req_index] <= req_tag;
          if (mem_add_read == 2'd3) begin
            valid[req_index][0] <= 1'b1;
            lru[req_index] <= 1'b1;  //way 0 was just used, so way 1 is LRU
          end

        //second line is empty
        end else if (~valid[req_index][1]) begin
          datas1[req_index][mem_add_read] <= i_mem_rdata;
          tags1[req_index] <= req_tag;
          if (mem_add_read == 2'd3) begin
            valid[req_index][1] <= 1'b1;
            lru[req_index] <= 1'b0;  //way 1 was just used, so way 0 is LRU
          end
        
        //neither are empty, evict lru
        end else begin
          if (lru[req_index] == 1'b0) begin
            datas0[req_index][mem_add_read] <= i_mem_rdata;
            tags0[req_index] <= req_tag;
            if (mem_add_read == 2'd3) begin
              lru[req_index] <= 1'b1;  //way 0 was just used, so way 1 is LRU
            end

          end else begin
            datas1[req_index][mem_add_read] <= i_mem_rdata;
            tags1[req_index] <= req_tag;
            if (mem_add_read == 2'd3) begin
              lru[req_index] <= 1'b0;  //way 1 was just used, so way 0 is LRU
            end

          end
        end

        mem_add_read <= mem_add_read + 1;
      end
    end
  end


  //write signal to be set to 1 inside the state machine when in the write
  //state
  always @(*) begin
    //default values
    next_state = state;
    busy1 = 1'b0;
    case (state)
      IDLE: begin
        //if the CPU requests a write (i_req_wen) or a read (i_req_ren), AND
        //it doesn't hit, then needs to read from the main memory
        //NOTE: to read 4 sequential adresses in memory, needs a seperate
        //state?
        //might be easier if there are additional states
        if ((i_req_wen || i_req_ren) && ~hit) begin
          next_state = MEMREAD;
          busy1 = 1'b1;
        end

        //if write and hit, skip loading block into memory, go directly to
        //writing to both memory and cache
        if (hit && i_req_wen) begin
          next_state = MEMWRITE;
          busy1 = 1'b1;
        end
      end
      MEMREAD: begin
        //stay in memread as long as i_mem_ready is false?
        //NOTE: once you've read the final line (i.e, mem_add_read becomes
        //3 or 4 depending on indexing method, then transition to the next
        //state; you've finished reading the 4 blocks of data you need into
        //the cache)
        //
        //should transition out of MEMREAD once 4 words of data have been read
        //from the memory to the cache: i.e, once mem_add_read has reached
        //3 (or 4?)...
        //CASE i_req_ren_ff; during the request, it was simply a read; can
        //transition back to the idle state?
        //CASE i_req_wen_ff; recall that for a write
        //a) if miss, load block into memory, then write to both cache and
        //memory
        //b) if hit, write to both cache and memory. tbh idk how this would
        //really work
        busy1 = 1'b1;
        //after mem_add_read reaches 3, then should transition to next state
        //add
        //add+1
        //add+2
        //add+3
        if (mem_add_read == 3'd3) begin
          //once reading 4 words of data into the cache, if the initial
          //request was a read, transition back to idle state?
          if (i_req_ren_ff) begin
            next_state = IDLE;
            //otherwise, if the initial request was a write, then transition
            //to MEMWRITE state to write to both cache and memory?
          end else if (i_req_wen_ff) begin
            next_state = MEMWRITE;
          end
          busy1 = 1'b1;
        end
      end

      MEMWRITE: begin
        busy1 = 1'b1;
      end
    endcase
  end
endmodule

`default_nettype wire
//are request signals only present for one clk cycle ? 

//IDLE  --> MEMREAD --> 

//IDLE check request if hit complete in 1 cycle (read and write)
//Complete write through in one also? what if mem not ready ? 

//if not a hit always read memory (new state) (done for read)

//for write need to write back to memory 3rd state ? 
